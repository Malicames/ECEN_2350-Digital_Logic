`timescale 1ns / 1ps

//This is my top level and main module
module Main(
    input  clk,                     //Normal clock
    input  [4:0] btn,               //btn[0] resets everything
    input  [15:0] sw,               //sw[0] = P2, sw[15] = P1 
    output [15:0] led,              //LED array also used to display the game

    //7-segment display ports
    output [3:0] D0_AN,
    output [3:0] D1_AN,
    output [7:0] D0_SEG,
    output [7:0] D1_SEG,

    //HDMI stuff from the downloaded IP
    output hdmi_clk_n,              //Negative differential clock signal
    output hdmi_clk_p,              //Positive differential clock signal
    output [2:0] hdmi_tx_n,         //Negative transmission signal output
    output [2:0] hdmi_tx_p          //Positive Transmission signal output
);

    wire rst = btn[0];              //Button that is used to reset everything 
    wire clk_25MHz, clk_125MHz;     //25MHz for VGA signal and 125MHz for HDMI signal
    wire locked;                    //Locks the signal transmission until signal is stable
    wire sclk;                      //This is a slower clock for refreshing the screen animations
    wire hsync, vsync, vde;         //These wires carry output from vga_driver to input of hdmi converter
    wire [9:0] x_wire, y_wire;      //X and Y wires for general connections
    wire [7:0] R, G, B;             //Red, green, and blue signal that is carried to the input of HDMI converter
    wire game_over;                 //Game over signal from tug_of_war module

    //Clock wizard stuff
    clk_wiz_0 clkgen_inst (
        .clk_out1(clk_25MHz),       // 25 MHz pixel clock
        .clk_out2(clk_125MHz),      // 125 MHz for HDMI serializer
        .reset(rst),
        .locked(locked),
        .clk_in1(clk)
    );

    //Slower clock for the game display (100Hz)
    Clock100Hz slowclock (.clk(clk), .sclk(sclk));

    //Instances for the VGA driver module: Produces x,y in visible range
    vga_driver vga1 (
        .sysClock(clk),
        .clock25(clk_25MHz),
        .reset(rst),
        .hsync(hsync),
        .vsync(vsync),
        .vde(vde),
        .x(x_wire),
        .y(y_wire)
    );

    //Instances for tug_of_war module
    wire [3:0] flag_out;
    First game_first (
        .clk(clk),
        .sclk(sclk),
        .sw(sw),
        .btn(btn),
        .led(led),

        //7-Segment display ports through to the main module
        .D0_AN(D0_AN),
        .D1_AN(D1_AN),
        .D0_SEG(D0_SEG),
        .D1_SEG(D1_SEG),

        //Export flag and game_over
        .flag_out(flag_out),
        .game_over(game_over)
    );

    //Map flag_out (0..15) to screen X coordinate (flag center)
    localparam integer MIN_CENTER = 10'd45;      //Left-most flag center
    localparam integer MAX_CENTER = 10'd570;     //Right-most flag center

    //This ensures the flag is in the "center" at the beginning of every round
    wire [9:0] flag_center_x;
    assign flag_center_x = MIN_CENTER + ((flag_out * 10'd570) / 10'd15);

    //Image creator: renders checkerboards, rope, and triangle centered at flag_center_x
    image_creator (
        .clk(clk_25MHz),
        .sclk(sclk),
        .reset(rst),
        .game_over(game_over),
        .x(x_wire),
        .y(y_wire),
        .flag_center_x(flag_center_x),
        .red(R),
        .green(G),
        .blue(B)
    );

    //Instance for the VGA to HDMI converter module (the module is defined by the downloaded IP)
    hdmi_tx_0 Conversion (
      .pix_clk(clk_25MHz),      //Input wire from clock wizard
      .pix_clkx5(clk_125MHz),   //Input wire from clock wizard
      .pix_clk_locked(locked),  //Input wire that locks signal transmission until signal is stable
      .rst(rst),                //Reset input wire from main module input
      .red(R),                  //Input wire [7:0] R
      .green(G),                //Input wire [7:0] G
      .blue(B),                 //Input wire [7:0] B
      .hsync(hsync),            //Input wire hsync which is generated by the VGA driver
      .vsync(vsync),            //Input wire vsync which is generated by the VGA driver
      .vde(vde),                //Input wire vde which is generated by the VGA driver
      //.aux0_din(8'b0),          //Input wire [7:0] aux0_din which we will ignore since we don't have audio
      //.aux1_din(8'b0),          //Input wire [7:0] aux1_din which we will ignore since we don't have audio
      //.aux2_din(8'b0),          //Input wire [7:0] aux2_din which we will ignore since we don't have audio
      //.ade(1'b0),               //Input wire for audio data enable which we won't be using
      .TMDS_CLK_P(hdmi_clk_p),  //Outputs continuous square wave that acts as timing reference for the HDMI receiver (positive)
      .TMDS_CLK_N(hdmi_clk_n),  //Outputs continuous square wave that acts as timing reference for the HDMI receiver (negative)
      .TMDS_DATA_P(hdmi_tx_p),  //Output wire [2:0] TMDS_DATA_P this is pin hdmi_tx_p on the Boolean Board
      .TMDS_DATA_N(hdmi_tx_n)   //Output wire [2:0] TMDS_DATA_N this is pin hdmi_tx_n on the Boolean Board
    );

endmodule


//Passes flag_out and game_over up
module First(
    input clk,
    input sclk,
    input [15:0] sw,
    input [4:0] btn,
    output [15:0] led,

    output [3:0] D0_AN,
    output [3:0] D1_AN,
    output [7:0] D0_SEG,
    output [7:0] D1_SEG,

    output [3:0] flag_out,
    output game_over
);

    wire [15:0] flip_p1;
    wire [15:0] flip_p2;
    wire [3:0] flag_internal;
    wire game_over_internal;

    //Tug_of_war instances 
    tug_of_war (
        .clk(clk),
        .sclk(sclk),
        .btn_reset(btn[0]),
        .sw_p1(sw[0]),
        .sw_p2(sw[15]),
        .led(led),
        .flip_p1(flip_p1),
        .flip_p2(flip_p2),
        .flag_out(flag_internal),
        .game_over(game_over_internal),
        .D0_AN(D0_AN),
        .D1_AN(D1_AN),
        .D0_SEG(D0_SEG),
        .D1_SEG(D1_SEG)
    );

    assign flag_out = flag_internal;
    assign game_over = game_over_internal;

endmodule


//Tug_of_war (Runs on sclk and outputs flag_out and game_over)
module tug_of_war (
    input  wire        clk,
    input  wire        sclk,
    input  wire        btn_reset,
    input  wire        sw_p1,
    input  wire        sw_p2,

    output reg [15:0]  led,
    output reg [15:0]  flip_p1,
    output reg [15:0]  flip_p2,

    output reg          game_over,     //Outputs game_over (Had issues with this)
    output reg [3:0]    flag_out,      //Outputs flag position (Had issues with this)

    output [3:0] D0_AN,
    output [3:0] D1_AN,
    output [7:0] D0_SEG,
    output [7:0] D1_SEG
);

    //Game state
    reg [3:0] flag = 4'd8;

    reg sw_p1_prev = 0;
    reg sw_p2_prev = 0;

    reg [1:0] winner = 2'b00;

    //Initialize outputs
    initial begin
        flip_p1 = 16'b0;
        flip_p2 = 16'b0;
        led = 16'b0;
        flag_out = 4'd8;
        game_over = 1'b0;
        winner = 2'b00;
    end

    //Movement of triangle, switch flip counting, and win detection
    always @(posedge sclk or posedge btn_reset) begin
        if (btn_reset) begin
            flag      <= 4'd8;
            flip_p1   <= 16'd0;
            flip_p2   <= 16'd0;
            sw_p1_prev <= sw_p1;
            sw_p2_prev <= sw_p2;
            game_over <= 1'b0;
            winner    <= 2'b0;
        end else begin
            if (!game_over) begin
                //Player 1 switch flip counting using Edge detection
                if (sw_p1 != sw_p1_prev) begin
                    flip_p1 <= flip_p1 + 1;
                    if (flag > 0)
                        flag <= flag + 1;
                end

                //Player 2 switch flip counting also using edge detection
                if (sw_p2 != sw_p2_prev) begin
                    flip_p2 <= flip_p2 + 1;
                    if (flag < 15)
                        flag <= flag - 1;
                end

                //Update previous switch state
                sw_p1_prev <= sw_p1;
                sw_p2_prev <= sw_p2;

                //Win detection
                if (flag == 0) begin
                    game_over <= 1'b1;
                    winner <= 2'b01;
                end else if (flag == 15) begin
                    game_over <= 1'b1;
                    winner <= 2'b10;
                end
            end
        end
    end

    //LED display of flag position
    always @(*) begin
        led = 16'b0;
        led[15 - flag] = 1'b1;
    end

    //Outputs flag to flag_out synchronized to sclk
    always @(posedge sclk or posedge btn_reset) begin
        if (btn_reset) flag_out <= 4'd8;
        else flag_out <= flag;
    end

    //7-Segmnet display
    localparam [7:0] SEG_BLANK = 8'b11111111;
    localparam [7:0] SEG_1     = 8'b11111001;  
    localparam [7:0] SEG_2     = 8'b10100100;

    reg [7:0] seg_data;

    //Win celebration 
    always @(*) begin
        if (game_over) begin
            case (winner)
                2'b01: seg_data = SEG_1; //Player 1 wins
                2'b10: seg_data = SEG_2; //Player 2 wins
                default: seg_data = SEG_BLANK;
            endcase
        end else begin
            seg_data = SEG_BLANK; //Blank/off during gameplay
        end
    end

    //Enable all digits
    assign D0_AN = 8'b00000000;
    assign D1_AN = 8'b00000000;

    //Drive segment lines
    assign D0_SEG = seg_data;
    assign D1_SEG = seg_data;

endmodule

//This is what creates all the fun shapes as well as controls what the shapes do (partially)
module image_creator(
    input clk,          
    input sclk,        
    input reset,
    input game_over,           //Connects everything
    input [9:0] x,
    input [9:0] y,
    input [9:0] flag_center_x, 
    output reg [7:0] red,
    output reg [7:0] green,
    output reg [7:0] blue
    );

    //Triangle: Tells it to stop short of generating pixels as it goes down the triangle 
    localparam integer TRI_HALF_MAX = 25;
    localparam integer TRI_HEIGHT   = 50;

    localparam integer TRI_Y_TOP    = 225;
    localparam integer TRI_Y_BOTTOM = TRI_Y_TOP + TRI_HEIGHT;

    //Increments the flag down to zero
    integer dy;
    integer current_half;

    localparam integer LEFT_CB_END  = 48;
    localparam integer RIGHT_CB_BEG = 660 - 48;

    //Blink Registers for game over
    reg [23:0] blink_counter = 0;
    reg blink_on = 1'b1;

    always @(posedge clk) begin
        
        //If game is over begin blinking the flag if the blink is on
        if (game_over) begin
            blink_counter <= blink_counter + 1;
            //Toggle every 0.5s at 25MHz
            if (blink_counter >= 24'd12500000) begin
                blink_counter <= 0;
                blink_on <= ~blink_on;
            end
        end else begin
            blink_counter <= 0;
            blink_on <= 1'b1;
        end

        //Default Background
        red   <= 8'b00000000;
        green <= 8'b00000000;
        blue  <= 8'b00000000;

        //Left checkerboard (~16x16 tiles)
        //If the current pixel is in the left region of the screen
        //Then XOR every 4 pixels up and down
        //If we have XORed, begin making checker board pattern passed on XOR output
        //**We must always have 1 so we keep the least significant bit**
        if (x < LEFT_CB_END) begin
            if (((x >> 4) ^ (y >> 4)) & 1) begin
                red   <= 8'b11111111; green <= 8'b11111111; blue <= 8'b11111111;
            end else begin
                red   <= 8'b00000000; green <= 8'b00000000; blue <= 8'b00000000;
            end
        end

        //Right checkerboard (~16x16 tiles)
        else if (x >= RIGHT_CB_BEG && x < 660) begin
            if (((x >> 4) ^ (y >> 4)) & 1) begin
                red   <= 8'b11111111; green <= 8'b11111111; blue <= 8'b11111111;
            end else begin
                red   <= 8'b00000000; green <= 8'b00000000; blue <= 8'b00000000;
            end
        end

        //The rope
        else if (y >= 215 && y <= 225) begin
            red   <= 8'b11000000;   //210
            green <= 8'b10100000;   //180
            blue  <= 8'b10000000;   //140
        end

        //Calls the blinking functions and applies it when game_over = 1
        //Checks if the pixel row is inside the triangles vertical area 
        else if (y >= TRI_Y_TOP && y <= TRI_Y_BOTTOM) begin
            dy = y - TRI_Y_TOP; 
            //Computes how wide the triangle should be on that row 
            current_half = TRI_HALF_MAX - (dy * TRI_HALF_MAX) / TRI_HEIGHT;
 
            //Checks if the pixel column is inside the specified width 
            //Draws a red pixel only if the game is not over or if the game is over and the blink is on
            if ((!game_over || blink_on) &&
                x >= (flag_center_x - current_half) &&
                x <= (flag_center_x + current_half)) begin
                red   <= 8'b11111111;
                green <= 8'b00000000;
                blue  <= 8'b00000000;
            end
        end
    end
endmodule

//VGA driver for the HDMI stuff
module vga_driver (
    input wire sysClock,
    input wire clock25,   //25Mhz
    input wire reset,     //Active high
    output reg vde,       //Video enable 
    output reg hsync,     //Horizontal sync 
    output reg vsync,     //Vertical sync
    output reg [9:0] x,y  //Position of pixels: x 0-799 and y 0-524 (for 480p)
     );

     //VGA timing values for 660x480 visible region
     parameter hor_display = 660;       //Pixels actually displayed
     parameter hor_fPorch = 48;         //Horizontal front porch (no pixels left of display)
     parameter hor_bPorch = 16;         //Horizontal back porch (no pixels right of display)
     parameter hor_retrace = 96;        //Horizontal retrace (cathode ray takes time to move)
     parameter hor_MAX = hor_display + hor_fPorch + hor_bPorch + hor_retrace - 1; //Max value of hoirzontal counter 799

     //Values for vertical display (525 pixels total)
     parameter ver_display = 480;       //Pixels actually displayed
     parameter ver_fPorch = 10;         //Vertical front porch (no pixels above display)
     parameter ver_bPorch = 33;         //Vertical front porch (no pixels below display)
     parameter ver_retrace = 2;         //Vertical retrace (cathode ray takes time to move)
     parameter ver_MAX = ver_display + ver_fPorch + ver_bPorch + ver_retrace - 1; //Max value of hoirzontal counter 524

     reg [9:0] h_count_reg = 0, h_count_next = 0;   //10 bits to for max value
     reg [9:0] v_count_reg = 0, v_count_next = 0;   //10 bits to for max value

     //Horizontal counter
     always @(posedge clock25 or posedge reset) begin
         if (reset) begin
             h_count_reg <= 0;
         end else begin
             if (h_count_reg == hor_MAX)
                 h_count_reg <= 0;
             else
                 h_count_reg <= h_count_reg + 1;
         end
     end

     //Vertical counter
     always @(posedge clock25 or posedge reset) begin
         if (reset) begin
             v_count_reg <= 0;
         end else begin
             if (h_count_reg == hor_MAX) begin
                 if (v_count_reg == ver_MAX)
                     v_count_reg <= 0;
                 else
                     v_count_reg <= v_count_reg + 1;
             end
         end
     end

     //This times the HDMI and VGA output making sure everything is synced
     //Uses the horizontal position to create hsync pulses
     //Uses the vertical position to create vsync pulses
     //Creates vde that is true when video pixels should be displayed
     //Shows the current pixel position on the X and Y axies 
     always @(*) begin
         hsync = (h_count_reg >= (hor_display + hor_bPorch) && h_count_reg <= (hor_display + hor_bPorch + hor_retrace - 1));
         vsync = (v_count_reg >= (ver_display + ver_bPorch) && v_count_reg <= (ver_display + ver_bPorch + ver_retrace - 1));
         vde   = (h_count_reg < hor_display) && (v_count_reg < ver_display);
         x = h_count_reg;
         y = v_count_reg;
     end

endmodule


//Slowclock100Hz: derive 100Hz from system clock
module Clock100Hz (input clk, output sclk);
    reg [31:0] counter = 0;
    reg hundredhertz = 1'b0;

    always @(posedge clk) begin
        counter <= counter + 1;
        if (counter >= 250000) begin
            counter <= 0;
            hundredhertz <= ~hundredhertz;
        end
    end

    assign sclk = hundredhertz;
endmodule
